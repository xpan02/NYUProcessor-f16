
----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    17:14:53 10/22/2016 
-- Design Name: 
-- Module Name:    InstructionMemory - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.std_logic_unsigned.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity InstructionMemory is
port(
     skey: in std_logic_vector(127 downto 0);
	  din: in std_logic_vector(63 downto 0);
     address: in std_logic_vector(31 downto 0);
	  Instruction: out std_logic_vector(31 downto 0));
	  
end InstructionMemory;
--IMM1=skey(31 downto 16)
--IMM2=skey(15 downto 0)
--IMM3=skey(63 downto 48)
--IMM4=skey(47 downto 32)
--IMM5=skey(95 downto 80)
--IMM6=skey(79 downto 64)
--IMM7=skey(127 downto 112)
--IMM8=skey(111 downto 96)
--offset1=L(0)DM(26)
--offset2=L(1)DM(27)
--offset3=L(2)Dm(28)
--offset4=L(3)DM(29)

architecture Behavioral of InstructionMemory is

type ramtype3 is array(0 to 171)of std_logic_vector(31 downto 0);
signal imem: ramtype3:=
(
 "00000000000000000000100000010000",--0 ADD RO,RO, R1 R1=0
 "00000000000000000001000000010000",--1 ADD R0,RO, R2 R2=0
 "00000000000000000001100000010000",--2 ADD RO,RO, R3 R3=0
 "00000100000111100000000000000000",--3 ****ADDI,RO,R30,skey(31 downto 16) R30=00..skey(31 downto 16)
 "00010111110111100000000000010000",--4 SHL R30 R30 16 R30=skey(31 downto 16)...000
 "00000100000111010000000000000000",--5 ****ADDI,RO,R29,SKEY(15 downto 0) R29=000.....skey(15 downto 0)
 "00000011110111011111000000010000",--6 ADD,R30 R29,R30 R30=skey(31 downto 0) 
 "00100000000111100000000000011010",--7 SW RO, R30 offset M[0+offset1]<-R30
 "00000100000111100000000000000000",--8 *****ADDI,RO,R30,skey(63 downto 48) R30=00..skey(63 downto 48)
 "00010111110111100000000000010000",--9 SHL R30 R30 16 R30=skey(63 downto 48)...000
 "00000100000111010000000000000000",--10 **** ADDI,RO,R29,SKEY(47 downto 32) R29=000.....skey(47 downto 32)
 "00000011110111011111000000010000",--11 ADD,R30 R29,R30 R30=skey(63 downto 32) 
 "00100000000111100000000000011011",--12 SW RO, R30 offset M[0+offset2]<-R30
 "00000100000111100000000000000000",--13 ****ADDI,RO,R30,skey(95 downto 80) R30=00..skey(95 downto 80)
 "00010111110111100000000000010000",--14 SHL R30 R30 16 R30=skey(95 downto 80)...000
 "00000100000111010000000000000000",--15 **** ADDI,RO,R29,SKEY(79 downto 64) R29=000.....skey(79 downto 64)
 "00000011110111011111000000010000",--16 ADD,R30 R29,R30 R30=skey(95 downto 64) 
 "00100000000111100000000000011100",--17 SW RO, R30 offset M[0+offset3]<-R30
 "00000100000111100000000000000000",--18 ******ADDI,RO,R30,skey(127 downto 112) R30=00..skey(127 downto 112)
 "00010111110111100000000000010000",--19 SHL R30 R30 16 R30=skey(127 downto 112)...000
 "00000100000111010000000000000000",--20******* ADDI,RO,R29,SKEY(111 downto 96) R29=000.....skey(111 downto 96)
 "00000011110111011111000000010000",--21 ADD,R30 R29,R30 R30=skey(127 downto 96) 
 "00100000000111100000000000011101",--22 SW RO, R30 offset M[0+offset4]<-R30
 "00000100000101010000000000000100",--23 ADDI,RO,R21,4 R21=4
 "00000100000101100000000000011010",--24 ADDI RO R22,26 R22=26
 "00000100000101110000000001001110",--25 ADDI R0 R23,78 R23=78
 "00000000000000000010000000010000",--26 ADD RO RO R4 R4=0
 "00000000000000000010100000010000",--27 ADD RO RO R5 R5=0
 "00011100010010000000000000000000",--28 R8<-MEM[R2+IMM_S)
 "00011100001010010000000000011010",--29 R9<-MEM(R1+IMM_l)
 "00000000100001010011000000010000",--30 ADD R4 R5,R6
 "00000001000001100101000000010000",--31 ADD R8 R6 R10
 "00000100000010110000000000000011",--32 ADDI RO R11 3
 "00000000000000000110000000010000",--33 ADD RO RO R12
 "00101001011011000000000000000101",--34 BEQ R11 R12 IMM
 "00010101010011010000000000000001",--35 SHL R10 R31 1
 "00011001010011100000000000011111",--36 SHR R10 R13 1
 "00000001101011100101000000010000",--37 ADD R13 R14 31
 "00000101100011000000000000000001",--38 ADDI R12 R12 1
 "00110000000000000000000000100010",--39 JMP IMM
 "00100000010010100000000000000000",--40 SW R2 R10 IMM_S branch here
 "00000000000010100010000000010000",--41 add RO R10 R4
 "00000000100001010011000000010000",--42 add R4 R5 R6
 "00000001001001100101000000010000",--43 add R9 R6 R10
 "00001100110010110000000000011111",--44 ANDI R6 R11 00....11111
 "00000000000000000110000000010000",--45 AND RO RO R12
 "00101001011011000000000000000101",--46 bEQ R11 R12 IMM
 "00010101010011010000000000000001",--47 SHL R10 R13 1
 "00011001010011100000000000011111",--48 SHR R10 R14 31
 "00000001101011100101000000010000",--49 ADD R13 R14 R10
 "00000101100011000000000000000001",--50 ADDI R12 R12 1
 "00110000000000000000000000101110",--51 JMP IMM
 "00100000001010100000000000011010",--52 SW R1 R10 IMML branch here
 "00000000000010100010100000010000",--53 ADD RO R10 R5
 "00000100001000010000000000000001",--54 ADDI R1 R1 1
 "00000100010000100000000000000001",--55 ADDI R2 R2 1
 "00000100011000110000000000000001",--56 ADDI R3 R3 1
 "00101100001101010000000000000001",--57 BNE R1 R21 IMM
 "00000000000000000000100000010000",--58 ADD RO RO R1
 "00101100010101100000000000000001",--59 BNE R2 R22 IMM
 "00000000000000000001000000010000",--60 ADD RO RO R2
 "00101000011101110000000000000001",--61 BEQ R3 R22 IMM
 "00110000000000000000000000011100",--62 JMP RETURN
 "00000000000000000001100000010000",--63 ADD RO RO R3
  -- end of key expension start of RC5-enc
 "00000100000111100000000000011010",--64 ADDI R0 R30 26 R30=26
 "00000000000000000010000000010000",--65 ADD RO RO R4 R4=0
 "00000000000000000010100000010000",--66 ADD RO RO R5 R5=0
 "00000100000001000000000000000000",--67 addi RO R4 din(63 downto 48)
 "00010100100001000000000000010000",--68 SHL R4 R4 16
 "00000100000111010000000000000000",--69 ADDI RO R29 din(47 downto 32)
 "00000000100111010010000000010000",--70 add R4 R29,R4 r4=din(63 downto 32)
 "00000100000001010000000000000000",--71 addi RO R5 din(31 downto 16)
 "00010100101001010000000000010000",--72 SHL R5 R5 16
 "00000100000111010000000000000000",--73 ADDI RO R29 din(15 downto 0)
 "00000000101111010010100000010000",--74 add R5 R29,R5 r5=din(31 downto 0)
 "00011100011111110000000000000000",--75 lw r3 r31 offset r31=M[0+offset]
 "00000000100111110010000000010000",--76 ADD R4 R31 R4 r4=din(63 downto 32)+M[0+offset]
 "00011100011111110000000000000001",--77 LW R3 R31 OFFSET+1 R31=M[0 +offset+1]
 "00000000101111110010100000010000",--78 ADD R5 R31 R5 r5=din(31 downto 0)+M[0+offset+1]
 "00000100011000110000000000000010",--79 addi r3 r3 2,r3=2
 "00000000100000000011000000010100",--80 NOR R4 RO R6  //RETURN
 "00000000101000000011100000010100",--81 NOR R5 RO R7
 "00000000100001110011100000010010",--82 ADD R4 R7 R7
 "00000000101001100011000000010010",--83 AND R5 R6 R6
 "00000000110001110100000000010000",--84 ADD R6 R7 R8 R8==AB_XOR
 "00001100101001110000000000011111",--85 ANDI R5 R7 000..111
 "00000000000000000011000000010000",--86 ADD RO RO R6
 "00000000000010000100100000010000",--87 ADD RO R8 R9
 "00101000110001110000000000000101",--88 BEQ R6 R7 IMM JUMP HERE
 "00010101001010100000000000000001",--89 SHL R9 R10 1
 "00011001001010110000000000011111",--90 SHR R9 R11 31
 "00000001010010110100100000010000",--91 ADD R10 R11 R9
 "00000100110001100000000000000001",--92 ADDI R6 R6 1
 "00110000000000000000000001011000",--93 JMP 88
 "00011100011111110000000000000000",--94 LW R3 R31 OFFSET
 "00000001001111110010000000010000",--95 ADD R9 R31 R4
 "00000000100000000011000000010100",--96 NOR R4 RO R6
 "00000000101000000011100000010100",--97 nor r5 ro r7
 "00000000100001110011100000010010",--98 aNd r4 r7 r7
 "00000000101001100011000000010010",--99 aNd r5 r6 r6
 "00000000110001110110000000010000",--100 ADD R6 R7 R12
 "00001100100001110000000000011111",--101 ANDI R4 R7 000..11111
 "00000000000000000011000000010000",--102 ADD RO RO R6
 "00000000000011000110100000010000",--103 ADD RO R12 R13
 "00101000110001110000000000000101",--104 BRANCH
 "00010101101010100000000000000001",--105 SHL R13 R10 1
 "00011001101010110000000000011111",--106 SHR R13 R11 31
 "00000001010010110110100000010000",--107 ADD R1O R11 R13
 "00000100110001100000000000000001",--108 ADDI R6 R6 1
 "00110000000000000000000001101000",--109 JUMP TO BEANCH 104
 "00011100011111110000000000000001",--110 lW R3 R31 OFFSET+1
 "00000001101111110010100000010000",--111 ADD R13 R31 R5
 "00000100011000110000000000000010",--112 ADDI R3 R3 2
 "00101000011111100000000000000001",--113 BEQ 115
 "00110000000000000000000001010000",--114 JUMP 80
 "00000000000000001000100000010000",--115 R17=0
 "00000000000000001001000000010000",--116 R18=0
 "00000000000001001000100000010000",--117 R17 store the final result of A
 "00000000000001011001000000010000",--118 R18 store the final result of B
 -- end of encrtpyion start of decryption
 "00000000000000000010000000010000",--119 add RO RO R4
 "00000000000000000010100000010000",--120 ADD RO RO R5
 "00000100000001000000000000000000",--121 addi RO R4 din(63 downto 48)
 "00010100100001000000000000010000",--122 SHL R4 R4 16
 "00000100000111010000000000000000",--123 ADDI RO R29 din(47 downto 32)
 "00000000100111010010000000010000",--124 add R4 R29,R4 r4=din(63 downto 32)
 "00000100000001010000000000000000",--125 addi RO R5 din(31 downto 16)
 "00010100101001010000000000010000",--126 SHL R5 R5 16
 "00000100000111010000000000000000",--127 ADDI RO R29 din(15 downto 0)
 "00000000101111010010100000010000",--128 add R5 R29,R5 r5=din(31 downto 0)
 "00000100000000110000000000011000",--129 ADDI RO R3 24
 "00011100011010000000000000000001",--130 LW R3 R8 OFFSET+1 R8<=S[25] RETURN
 "00000000101010000011100000010001",--131 SUB R5 R8 R7 R7=B-S[25]
 "00001100100010010000000000011111",--132 ANDI R4 R9 000...11111 R9 SHIFT BITS
 "00000000000000000100000000010000",--133 ADD RO RO R8 r8=0
 "00000000000001110101100000010000",--134 ADD RO R7 R11 R11=R7=B-s[25]
 "00101001000010010000000000000101",--135 BEQ R8 R9 IMM=5
 "00011001011011000000000000000001",--136 SHR R11 R12 1
 "00010101011011010000000000011111",--137 SHL R11 R13 31
 "00000001100011010101100000010000",--138 ADD R12 R13 R11
 "00000101000010000000000000000001",--139 ADDI R8 R8 1
 "00110000000000000000000010000111",--140 JMP 135
 "00000000100000000100000000010100",--141 NOR R4 R0 R8
 "00000001011000000100100000010100",--142 NOR R11 R0 R9
 "00000000100010010100100000010010",--143 AND R4 R9 R9
 "00000001000010110100000000010010",--144 AnD R8 R11 R8
 "00000001000010010010100000010000",--145 ADD R8 R9 R5
 "00011100011010000000000000000000",--145 LW R3 R8 OFFSET
 "00000000100010000011000000010001",--147 SUB R4 R8 R6 R6=a-s[24]
 "00001100101010010000000000011111",--148 ANDI R5 R9 000.11111 
 "00000000000000000100000000010000",--149 ADD RO RO R8
 "00000000000001100101000000010000",--150 ADD RO R6 R10
 "00101001000010010000000000000101",--151 BEQ R8 R9 5
 "00011001010011000000000000000001",--152 SHR R10 R12 1
 "00010101010011010000000000011111",--153 SHL R10 R13 31
 "00000001100011010101000000010000",--154 ADD R12 R13 R10 R10=(A-S[24]>>>B)
 "00000101000010000000000000000001",--155 ADDI R8 R8 1
 "00110000000000000000000010010111",--156 JUMP 151
 "00000001010000000100000000010100",--157 NOR R10 R0 R8
 "00000000101000000100100000010100",--158 NOR R5 R0 R9
 "00000001010010010100100000010010",--159 AND R10 R9 R9
 "00000000101010000100000000010010",--160 AND R5 R8 R8
 "00000001000010010010000000010000",--161 ADD R8 R9 R4
 "00001000011000110000000000000010",--162 SUBI R3 R3 2
 "00101000011000000000000000000001",--163 BEQ R3 R0 1
 "00110000000000000000000010000010",--164 JUMP RETURN 130
 "00011100011010000000000000000001",--165 LW R3 R8 OFFSET+1
 "00000000101010000010100000010001",--166 SUB R5 R8 R5
 "00011100011010000000000000000000",--167 LW R3 R8 OFFSET
 "00000000100010000010000000010001",--168 SUB R4 R8 R4
 "00000000000001011100100000010000",--169 ADD RO R5 R25 store dey result b in R[25]
 "00000000000001001100000000010000", --170 ADD RO R4 R24 store dey result A in R[24]
 "11111100000000000000000000000000" --171 halt
 );
 
begin
    imem(3)<="0000010000011110"&skey(31 downto 16);
	 imem(5)<="0000010000011101"&skey(15 downto 0);
	 imem(8)<="0000010000011110"&skey(63 downto 48);
	 imem(10)<="0000010000011101"&skey(47 downto 32);
	 imem(13)<="0000010000011110"&skey(95 downto 80);
	 imem(15)<="0000010000011101"&skey(79 downto 64);
	 imem(18)<="0000010000011110"&skey(127 downto 112);
	 imem(20)<="0000010000011101"&skey(111 downto 96);
	 imem(67)<="0000010000000100"&din(63 downto 48);
	 imem(69)<="0000010000011101"&din(47 downto 32);
	 imem(71)<="0000010000000101"&din(31 downto 16);
	 imem(73)<="0000010000011101"&din(15 downto 0);
	 imem(121)<="0000010000000100"&din(63 downto 48);
	 imem(123)<="0000010000011101"&din(47 downto 32);
	 imem(125)<="0000010000000101"&din(31 downto 16);
	 imem(127)<="0000010000011101"&din(15 downto 0);			 
    Instruction<=imem(conv_integer(address));

end Behavioral;